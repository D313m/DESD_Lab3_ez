library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use ieee.numeric_std.all;

entity moving_average_filter_en is
	generic (
		-- Filter order expressed as 2^(FILTER_ORDER_POWER)
		FILTER_ORDER_POWER : integer  := 5;
		TDATA_WIDTH        : positive := 24
	);
	Port (
		aclk          : in  std_logic;
		aresetn       : in  std_logic;
		
		s_axis_tvalid : in  std_logic;
		s_axis_tdata  : in  std_logic_vector(TDATA_WIDTH - 1 downto 0);
		s_axis_tlast  : in  std_logic;
		s_axis_tready : out std_logic;
		
		m_axis_tvalid : out std_logic;
		m_axis_tdata  : out std_logic_vector(TDATA_WIDTH - 1 downto 0);
		m_axis_tlast  : out std_logic;
		m_axis_tready : in  std_logic;
		
		enable_filter : in std_logic
	);
end moving_average_filter_en;

architecture Behavioral of moving_average_filter_en is
	component moving_average_filter is
		generic (
			-- Filter order expressed as 2^(FILTER_ORDER_POWER)
			FILTER_ORDER_POWER : integer  := 5;
			TDATA_WIDTH        : positive := 24
		);
		Port (
			aclk          : in  std_logic;
			aresetn       : in  std_logic;
			
			s_axis_tvalid : in  std_logic;
			s_axis_tdata  : in  std_logic_vector(TDATA_WIDTH - 1 downto 0);
			s_axis_tlast  : in  std_logic;
			s_axis_tready : out std_logic;
			
			m_axis_tvalid : out std_logic;
			m_axis_tdata  : out std_logic_vector(TDATA_WIDTH - 1 downto 0);
			m_axis_tlast  : out std_logic;
			m_axis_tready : in  std_logic
		);
	end component moving_average_filter;
	
	component all_pass_filter is
		generic (
			TDATA_WIDTH   : positive := 24
		);
		Port (
			aclk          : in  std_logic;
			aresetn       : in  std_logic;
			
			s_axis_tvalid : in  std_logic;
			s_axis_tdata  : in  std_logic_vector(TDATA_WIDTH - 1 downto 0);
			s_axis_tlast  : in  std_logic;
			s_axis_tready : out std_logic;
			
			m_axis_tvalid : out std_logic;
			m_axis_tdata  : out std_logic_vector(TDATA_WIDTH - 1 downto 0);
			m_axis_tlast  : out std_logic;
			m_axis_tready : in  std_logic
		);
	end component all_pass_filter;
	
begin
	
end Behavioral;